-- Stack Pointer Controller
